library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux_2_16 is
	Port(
			in0, in1 : in STD_LOGIC_VECTOR(15 downto 0);
			s : in STD_LOGIC;
			z : out STD_LOGIC_VECTOR(15 downto 0)
		);
end mux_2_16;

architecture Behavioral of mux_2_16 is

begin

	z <= 	in0 after 5ns when s = '0' else
			in1 after 5ns when s = '1' else
			x"0000" after 5ns;

end Behavioral;

